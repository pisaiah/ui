module iui

import gx

// Checkbox - implements Component interface
pub struct Switch {
	Component_A
pub mut:
	text     string
	bind_val &bool = unsafe { nil }
	cut      int   = 4
	thumb_x  int
}

pub fn (mut s Switch) get_thumb_x(g &GraphicsContext) int {
	if s.is_selected && s.thumb_x < s.height + s.cut {
		s.thumb_x += 2
		g.refresh_ui()
	}

	if !s.is_selected && s.thumb_x > s.cut {
		s.thumb_x -= 2
		g.refresh_ui()
	}

	return s.x + s.thumb_x
}

pub fn (mut s Switch) bind_to(val &bool) {
	unsafe {
		s.bind_val = val
	}
}

pub fn (mut s Switch) update_bind() {
	if isnil(s.bind_val) {
		return
	}

	unsafe {
		*s.bind_val = s.is_selected
	}
}

@[params]
pub struct SwitchConfig {
pub:
	bounds   Bounds
	selected bool
	text     string
}

pub fn Switch.new(cf SwitchConfig) &Switch {
	return &Switch{
		text:        cf.text
		x:           cf.bounds.x
		y:           cf.bounds.y
		width:       cf.bounds.width
		height:      cf.bounds.height
		is_selected: cf.selected
		thumb_x:     0
	}
}

// Get border color
fn (this &Switch) get_border(is_hover bool, ctx &GraphicsContext) gx.Color {
	if this.is_mouse_down {
		return ctx.theme.button_border_click
	}

	if is_hover {
		return ctx.theme.button_border_hover
	}
	return ctx.theme.button_border_normal
}

// Get background color
fn (this &Switch) get_background(is_hover bool, ctx &GraphicsContext) gx.Color {
	if this.is_selected {
		if this.is_mouse_down {
			return ctx.theme.accent_fill_third
		}
		if is_hover {
			return ctx.theme.accent_fill_second
		}
		return ctx.theme.accent_fill
	}

	if this.is_mouse_down {
		return ctx.theme.button_bg_click
	}

	if this.is_selected {
		return ctx.theme.accent_fill
	}

	if is_hover {
		return ctx.theme.button_bg_hover
	}

	return ctx.theme.button_bg_normal
}

// Draw Switch
pub fn (mut com Switch) draw(ctx &GraphicsContext) {
	// Draw Background & Border
	com.draw_background(ctx)

	// Detect click
	if com.is_mouse_rele {
		com.is_mouse_rele = false
		com.is_selected = !com.is_selected
		invoke_switch(com, ctx)
		com.update_bind()
	}

	if !isnil(com.bind_val) {
	}
	if !isnil(com.bind_val) {
		if com.is_selected != com.bind_val {
			com.is_selected = com.bind_val
		}
	}

	if com.thumb_x == 0 {
		com.thumb_x = if com.is_selected { com.height + com.cut } else { com.cut }
	}

	// Draw thumb/handle
	tx := com.get_thumb_x(ctx)
	wid := com.height - com.cut * 2
	ctx.gg.draw_rounded_rect_filled(tx, com.y + com.cut, wid, wid, 64, ctx.theme.button_border_normal)
	ctx.gg.draw_rounded_rect_filled(tx + 1, com.y + com.cut + 1, wid - 2, wid - 2, 64,
		ctx.theme.button_bg_normal)

	// Draw text
	com.draw_text(ctx)
}

// Draw background & border of Switch
fn (sw &Switch) draw_background(ctx &GraphicsContext) {
	is_hover := is_in(sw, ctx.win.mouse_x, ctx.win.mouse_y)

	bg := sw.get_background(is_hover, ctx)
	border := sw.get_border(is_hover, ctx)

	bh := sw.height * 2
	h := sw.height

	ctx.gg.draw_rounded_rect_filled(sw.x, sw.y, bh, h, 16, border)
	ctx.gg.draw_rounded_rect_filled(sw.x + 1, sw.y + 1, bh - 2, h - 2, 16, bg)
}

// Draw the text of Switch
fn (this &Switch) draw_text(ctx &GraphicsContext) {
	sizh := ctx.line_height / 2 // ctx.gg.text_height(this.text) / 2
	left := this.height * 2

	ctx.draw_text(this.x + left + 4, this.y + (this.height / 2) - sizh, this.text, ctx.font,
		gx.TextCfg{
		size:  ctx.font_size
		color: ctx.theme.text_color
	})
}

fn (sw &Switch) draw_circ(o int, g &GraphicsContext) {
}

pub struct SwitchEvent {
	ComponentEventGeneric[Switch]
}

pub fn invoke_switch(sw &Switch, ctx &GraphicsContext) {
	ev := SwitchEvent{
		target: sw
		ctx:    ctx
	}

	for f in sw.events.event_map['change'] {
		f(ev)
	}
}
