module file_dialog

#flag -I @VMODROOT/src/extra/file_dialog/

// TODO
pub fn color_picker() string {
	return ''
}

fn cstr(the_string string) &char {
	return &char(the_string.str)
}

// TODO
pub fn save_dialog(title string) string {
	return ''
}

// TODO
pub fn select_folder_dialog(title string, current string) string {
	return ''
}
