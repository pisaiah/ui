module extra

import iui as ui

struct Svg {
}