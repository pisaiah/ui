module iui

import gg

// Modal - implements Component interface
pub struct Modal {
	Component_A
pub mut:
	text       string
	needs_init bool
	close      &Button
	shown      bool
	close_idx  ?int

	in_width          int
	in_height         int
	left_off          int
	top_off           int = 50
	xs                int
	pack              bool
	container_pass_ev bool = true
	on_resize         ?fn (voidptr)
}

@[params]
pub struct ModalConfig {
pub:
	children  ?[]Component
	title     string
	width     int = 500
	height    int = 300
	left      int
	top       int = 50
	close_idx ?int
	on_resize ?fn (voidptr)
}

pub fn Modal.new(c ModalConfig) &Modal {
	return &Modal{
		text:       c.title
		z_index:    500
		needs_init: true
		in_width:   c.width
		in_height:  c.height
		close:      unsafe { nil }
		close_idx:  c.close_idx
		left_off:   c.left
		top_off:    c.top
		children:   c.children or { []Component{} }
		on_resize:  c.on_resize
	}
}

pub fn (mut this Modal) pack() {
	this.pack = true
}

pub fn (mut m Modal) calc_resize(ctx &GraphicsContext, ws gg.Size) {
	m.width = ws.width
	m.height = ws.height

	m.xs = (ws.width / 2) - (m.in_width / 2) - m.left_off
	if m.on_resize != none {
		mut ev := &DrawEvent{
			target: m
			ctx:    ctx
		}
		m.on_resize(ev)
	}
}

const modal_transparent = gg.rgba(0, 0, 0, 170)

pub fn (mut m Modal) draw(ctx &GraphicsContext) {
	ws := gg.window_size()

	if m.width != ws.width || m.height != ws.height {
		m.calc_resize(ctx, ws)
	}

	if m.z_index <= 501 {
		// Only draw background for one modal.
		ctx.gg.draw_rect_filled(0, 0, ws.width, ws.height, modal_transparent)
	}

	wid := m.in_width
	hei := m.in_height
	bord_wid := 5
	wid_2 := wid - (bord_wid * 2)
	bg := ctx.theme.textbox_border

	top := 28
	ctx.gg.draw_rounded_rect_filled(m.xs, m.top_off, wid, hei + bord_wid + top, 9, bg)

	ttop := m.top_off + (ctx.line_height / 2) - 1

	ctx.gg.draw_text(m.xs + 6, ttop, m.text, gg.TextCfg{
		size:  ctx.font_size
		color: ctx.theme.text_color
	})

	ctx.gg.draw_rect_filled(m.xs + bord_wid, m.top_off + top, wid_2, hei, ctx.theme.background)
	ctx.gg.draw_rect_empty(m.xs + bord_wid, m.top_off + top, wid_2, hei, ctx.theme.button_bg_click)

	mut app := ctx.win

	// Do component draw event again to fix z-index
	// if !isnil(m.draw_event_fn) {
	// m.draw_event_fn(mut app, &Component(m))
	// }

	if m.needs_init {
		if m.close_idx == none {
			m.make_close_btn(true)
		}
		m.needs_init = false
	}

	y_off := m.y + m.top_off + top
	for i, mut kid in m.children {
		kid.draw_event_fn(mut app, kid)
		kid.draw_with_offset(ctx, m.xs, y_off + 2)

		if m.pack {
			if kid.width > m.in_width {
				m.in_width = kid.width + (kid.x * 2)
				if !isnil(m.close) {
					m.close.x = m.in_width - 115
				} else if m.close_idx != none {
					if i == m.close_idx {
						kid.x = m.in_width - 115
					}
				}
				m.calc_resize(ctx, ws)
			}
		}
	}
}

pub fn (mut this Modal) make_close_btn(ce bool) &Button {
	mut close := Button.new(
		text:   'OK'
		bounds: Bounds{200, this.in_height - 40, 100, 30}
	)

	if 300 > this.in_width {
		close.x = this.in_width - 115
	}

	if ce {
		close.subscribe_event('mouse_up', default_modal_close_fn)
		if this.needs_init {
			close.is_action = true
		}
	}

	this.children << close
	this.close = close
	return close
}

pub fn default_modal_close_fn(mut e MouseEvent) {
	e.ctx.win.components = e.ctx.win.components.filter(mut it !is Modal)
}
